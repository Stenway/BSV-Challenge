Hello�🌎�����Test 𝄞